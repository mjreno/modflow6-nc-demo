netcdf csub_sk03a {
dimensions:
	LINELENGTH = 300 ;
	LENAUXNAME = 16 ;
	LENBOUNDNAME = 40 ;
	LENTIMESERIESNAME = 40 ;
	NPER = 2 ;
	NLAY = 3 ;
	NROW = 21 ;
	NCOL = 20 ;
	NCPL = 420 ;
	NCELLDIM = 3 ;
	dim_chd_0_maxbound = 42 ;
	dim_chd_0_niper = 1 ;
variables:
	int dis_nlay ;
		dis_nlay:_FillValue = -2147483647 ;
		dis_nlay:mf6_input = "DIS6:CSUB_SK03A/DIS/NLAY" ;
	int dis_nrow ;
		dis_nrow:_FillValue = -2147483647 ;
		dis_nrow:mf6_input = "DIS6:CSUB_SK03A/DIS/NROW" ;
	int dis_ncol ;
		dis_ncol:_FillValue = -2147483647 ;
		dis_ncol:mf6_input = "DIS6:CSUB_SK03A/DIS/NCOL" ;
	double dis_delr(NCOL) ;
		dis_delr:_FillValue = 3.e+30 ;
		dis_delr:mf6_input = "DIS6:CSUB_SK03A/DIS/DELR" ;
	double dis_delc(NROW) ;
		dis_delc:_FillValue = 3.e+30 ;
		dis_delc:mf6_input = "DIS6:CSUB_SK03A/DIS/DELC" ;
	double dis_top(NLAY, NROW, NCOL) ;
		dis_top:_FillValue = 3.e+30 ;
		dis_top:mf6_input = "DIS6:CSUB_SK03A/DIS/TOP" ;
	double dis_botm(NLAY, NROW, NCOL) ;
		dis_botm:_FillValue = 3.e+30 ;
		dis_botm:mf6_input = "DIS6:CSUB_SK03A/DIS/BOTM" ;
	double ic_strt(NLAY, NROW, NCOL) ;
		ic_strt:_FillValue = 3.e+30 ;
		ic_strt:mf6_input = "IC6:CSUB_SK03A/IC/STRT" ;
	int npf_save_flows ;
		npf_save_flows:_FillValue = -2147483647 ;
		npf_save_flows:mf6_input = "NPF6:CSUB_SK03A/NPF/SAVE_FLOWS" ;
	int npf_save_specific_discharge ;
		npf_save_specific_discharge:_FillValue = -2147483647 ;
		npf_save_specific_discharge:mf6_input = "NPF6:CSUB_SK03A/NPF/SAVE_SPECIFIC_DISCHARGE" ;
	int npf_icelltype(NLAY, NROW, NCOL) ;
		npf_icelltype:_FillValue = -2147483647 ;
		npf_icelltype:mf6_input = "NPF6:CSUB_SK03A/NPF/ICELLTYPE" ;
	double npf_k(NLAY, NROW, NCOL) ;
		npf_k:_FillValue = 3.e+30 ;
		npf_k:mf6_input = "NPF6:CSUB_SK03A/NPF/K" ;
	double npf_k33(NLAY, NROW, NCOL) ;
		npf_k33:_FillValue = 3.e+30 ;
		npf_k33:mf6_input = "NPF6:CSUB_SK03A/NPF/K33" ;
	char chd_0_ts_filerecord(LINELENGTH) ;
		chd_0_ts_filerecord:_Encoding = "ascii" ;
		chd_0_ts_filerecord:mf6_input = "CHD6:CSUB_SK03A/CHD_0/TS_FILERECORD" ;
	int chd_0_maxbound ;
		chd_0_maxbound:_FillValue = -2147483647 ;
		chd_0_maxbound:mf6_input = "CHD6:CSUB_SK03A/CHD_0/MAXBOUND" ;
	int chd_0_cellid(dim_chd_0_niper, dim_chd_0_maxbound, NCELLDIM) ;
		chd_0_cellid:_FillValue = -2147483647 ;
		chd_0_cellid:mf6_input = "CHD6:CSUB_SK03A/CHD_0/CELLID" ;
	double chd_0_head(dim_chd_0_niper, dim_chd_0_maxbound) ;
		chd_0_head:_FillValue = 3.e+30 ;
		chd_0_head:mf6_input = "CHD6:CSUB_SK03A/CHD_0/HEAD" ;
		chd_0_head:mf6_timeseries = "chd_0_head_ts" ;
	char chd_0_head_ts(dim_chd_0_niper, dim_chd_0_maxbound, LENTIMESERIESNAME) ;
		chd_0_head_ts:_Encoding = "ascii" ;
	int chd_0_iper(dim_chd_0_niper) ;
		chd_0_iper:_FillValue = -2147483647 ;
		chd_0_iper:mf6_input = "CHD6:CSUB_SK03A/CHD_0/IPER" ;

// global attributes:
		:description = "MODFLOW 6 NetCDF4 file prototype" ;
		:history = "Created Mon Jan 22 09:06:31 2024" ;
		:source = "mf6netcdf4.py" ;
		:mf6_modeltype = "GWF6" ;
		:mf6_modelname = "CSUB_SK03A" ;
		:Conventions = "CF-1.8" ;
data:

 dis_nlay = 3 ;

 dis_nrow = 21 ;

 dis_ncol = 20 ;

 dis_delr = 0.5, 0.6, 0.72, 0.864, 1.0368, 1.24416, 1.492992, 1.7915904, 
    2.14990848, 2.579890176, 3.0958682112, 3.71504185344, 4.458050224128, 
    5.3496602689536, 6.41959232274432, 7.70351078729318, 9.24421294475182, 
    11.0930555337022, 13.3116666404426, 15 ;

 dis_delc = 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 
    50, 50, 50, 50, 50 ;

 dis_top =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 dis_botm =
  -12.1921110945163, -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, -12.1921110945163,
  -12.1921110945163, -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, -12.1921110945163,
  -12.1921110945163, -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, -12.1921110945163,
  -12.1921110945163, -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, -12.1921110945163,
  -12.1921110945163, -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, -12.1921110945163,
  -12.1921110945163, -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, -12.1921110945163,
  -12.1921110945163, -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, -12.1921110945163,
  -12.1921110945163, -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, -12.1921110945163,
  -12.1921110945163, -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, -12.1921110945163,
  -12.1921110945163, -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, -12.1921110945163,
  -12.1921110945163, -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, -12.1921110945163,
  -12.1921110945163, -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, -12.1921110945163,
  -12.1921110945163, -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, -12.1921110945163,
  -12.1921110945163, -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, -12.1921110945163,
  -12.1921110945163, -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, -12.1921110945163,
  -12.1921110945163, -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, -12.1921110945163,
  -12.1921110945163, -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, -12.1921110945163,
  -12.1921110945163, -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, -12.1921110945163,
  -12.1921110945163, -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, -12.1921110945163,
  -12.1921110945163, -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, -12.1921110945163,
  -12.1921110945163, -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, 
    -12.1921110945163, -12.1921110945163, -12.1921110945163, -12.1921110945163,
  -21.3361944154035, -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, -21.3361944154035,
  -21.3361944154035, -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, -21.3361944154035,
  -21.3361944154035, -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, -21.3361944154035,
  -21.3361944154035, -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, -21.3361944154035,
  -21.3361944154035, -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, -21.3361944154035,
  -21.3361944154035, -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, -21.3361944154035,
  -21.3361944154035, -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, -21.3361944154035,
  -21.3361944154035, -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, -21.3361944154035,
  -21.3361944154035, -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, -21.3361944154035,
  -21.3361944154035, -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, -21.3361944154035,
  -21.3361944154035, -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, -21.3361944154035,
  -21.3361944154035, -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, -21.3361944154035,
  -21.3361944154035, -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, -21.3361944154035,
  -21.3361944154035, -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, -21.3361944154035,
  -21.3361944154035, -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, -21.3361944154035,
  -21.3361944154035, -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, -21.3361944154035,
  -21.3361944154035, -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, -21.3361944154035,
  -21.3361944154035, -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, -21.3361944154035,
  -21.3361944154035, -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, -21.3361944154035,
  -21.3361944154035, -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, -21.3361944154035,
  -21.3361944154035, -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, 
    -21.3361944154035, -21.3361944154035, -21.3361944154035, -21.3361944154035,
  -30.4802777362907, -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, -30.4802777362907,
  -30.4802777362907, -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, -30.4802777362907,
  -30.4802777362907, -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, -30.4802777362907,
  -30.4802777362907, -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, -30.4802777362907,
  -30.4802777362907, -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, -30.4802777362907,
  -30.4802777362907, -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, -30.4802777362907,
  -30.4802777362907, -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, -30.4802777362907,
  -30.4802777362907, -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, -30.4802777362907,
  -30.4802777362907, -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, -30.4802777362907,
  -30.4802777362907, -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, -30.4802777362907,
  -30.4802777362907, -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, -30.4802777362907,
  -30.4802777362907, -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, -30.4802777362907,
  -30.4802777362907, -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, -30.4802777362907,
  -30.4802777362907, -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, -30.4802777362907,
  -30.4802777362907, -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, -30.4802777362907,
  -30.4802777362907, -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, -30.4802777362907,
  -30.4802777362907, -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, -30.4802777362907,
  -30.4802777362907, -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, -30.4802777362907,
  -30.4802777362907, -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, -30.4802777362907,
  -30.4802777362907, -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, -30.4802777362907,
  -30.4802777362907, -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, 
    -30.4802777362907, -30.4802777362907, -30.4802777362907, -30.4802777362907 ;

 ic_strt =
  -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018,
  -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018,
  -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018,
  -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018,
  -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018,
  -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018,
  -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018,
  -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018,
  -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018,
  -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018,
  -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018,
  -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018,
  -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018,
  -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018,
  -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018,
  -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018,
  -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018,
  -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018,
  -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018,
  -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018,
  -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018,
  -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018,
  -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018,
  -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018,
  -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018,
  -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018,
  -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018,
  -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018,
  -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018,
  -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018,
  -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018,
  -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018,
  -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018,
  -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018,
  -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018,
  -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018,
  -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018,
  -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018,
  -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018,
  -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018,
  -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018,
  -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018,
  -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018,
  -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018,
  -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018,
  -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018,
  -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018,
  -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018,
  -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018,
  -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018,
  -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018,
  -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018,
  -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018,
  -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018,
  -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018,
  -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018,
  -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018,
  -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018,
  -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018,
  -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018,
  -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018,
  -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018,
  -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, 
    -10.6680972077018, -10.6680972077018, -10.6680972077018, -10.6680972077018 ;

 npf_save_flows = 1 ;

 npf_save_specific_discharge = 1 ;

 npf_icelltype =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 npf_k =
  1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05,
  1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05,
  1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05,
  1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05,
  1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05,
  1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05,
  1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05,
  1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05,
  1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05,
  1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05,
  1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05,
  1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05,
  1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05,
  1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05,
  1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05,
  1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05,
  1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05,
  1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05,
  1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05,
  1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05,
  1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05, 1.7639049615909e-05, 
    1.7639049615909e-05, 1.7639049615909e-05,
  3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09,
  3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09,
  3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09,
  3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09,
  3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09,
  3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09,
  3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09,
  3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09,
  3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09,
  3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09,
  3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09,
  3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09,
  3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09,
  3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09,
  3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09,
  3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09,
  3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09,
  3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09,
  3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09,
  3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09,
  3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09, 3.5278099231818e-09, 
    3.5278099231818e-09, 3.5278099231818e-09,
  5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05,
  5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05,
  5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05,
  5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05,
  5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05,
  5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05,
  5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05,
  5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05,
  5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05,
  5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05,
  5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05,
  5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05,
  5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05,
  5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05,
  5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05,
  5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05,
  5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05,
  5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05,
  5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05,
  5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05,
  5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05, 5.2917148847727e-05, 
    5.2917148847727e-05, 5.2917148847727e-05 ;

 npf_k33 =
  1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06,
  1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06,
  1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06,
  1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06,
  1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06,
  1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06,
  1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06,
  1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06,
  1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06,
  1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06,
  1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06,
  1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06,
  1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06,
  1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06,
  1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06,
  1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06,
  1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06,
  1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06,
  1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06,
  1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06,
  1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06, 1.7639049615909e-06, 
    1.7639049615909e-06, 1.7639049615909e-06,
  3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10,
  3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10,
  3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10,
  3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10,
  3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10,
  3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10,
  3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10,
  3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10,
  3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10,
  3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10,
  3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10,
  3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10,
  3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10,
  3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10,
  3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10,
  3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10,
  3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10,
  3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10,
  3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10,
  3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10,
  3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10, 3.5278099231818e-10, 
    3.5278099231818e-10, 3.5278099231818e-10,
  5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06,
  5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06,
  5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06,
  5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06,
  5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06,
  5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06,
  5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06,
  5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06,
  5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06,
  5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06,
  5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06,
  5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06,
  5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06,
  5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06,
  5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06,
  5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06,
  5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06,
  5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06,
  5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06,
  5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06,
  5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06, 5.2917148847727e-06, 
    5.2917148847727e-06, 5.2917148847727e-06 ;

 chd_0_ts_filerecord = "csub_sk03a.ch.ts                                                                                                                                                                                                                                                                                            " ;

 chd_0_maxbound = 42 ;

 chd_0_cellid =
  1, 1, 20,
  1, 2, 20,
  1, 3, 20,
  1, 4, 20,
  1, 5, 20,
  1, 6, 20,
  1, 7, 20,
  1, 8, 20,
  1, 9, 20,
  1, 10, 20,
  1, 11, 20,
  1, 12, 20,
  1, 13, 20,
  1, 14, 20,
  1, 15, 20,
  1, 16, 20,
  1, 17, 20,
  1, 18, 20,
  1, 19, 20,
  1, 20, 20,
  1, 21, 20,
  3, 1, 20,
  3, 2, 20,
  3, 3, 20,
  3, 4, 20,
  3, 5, 20,
  3, 6, 20,
  3, 7, 20,
  3, 8, 20,
  3, 9, 20,
  3, 10, 20,
  3, 11, 20,
  3, 12, 20,
  3, 13, 20,
  3, 14, 20,
  3, 15, 20,
  3, 16, 20,
  3, 17, 20,
  3, 18, 20,
  3, 19, 20,
  3, 20, 20,
  3, 21, 20 ;

 chd_0_head =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 chd_0_head_ts =
  "chd                                     ",
  "chd                                     ",
  "chd                                     ",
  "chd                                     ",
  "chd                                     ",
  "chd                                     ",
  "chd                                     ",
  "chd                                     ",
  "chd                                     ",
  "chd                                     ",
  "chd                                     ",
  "chd                                     ",
  "chd                                     ",
  "chd                                     ",
  "chd                                     ",
  "chd                                     ",
  "chd                                     ",
  "chd                                     ",
  "chd                                     ",
  "chd                                     ",
  "chd                                     ",
  "chd                                     ",
  "chd                                     ",
  "chd                                     ",
  "chd                                     ",
  "chd                                     ",
  "chd                                     ",
  "chd                                     ",
  "chd                                     ",
  "chd                                     ",
  "chd                                     ",
  "chd                                     ",
  "chd                                     ",
  "chd                                     ",
  "chd                                     ",
  "chd                                     ",
  "chd                                     ",
  "chd                                     ",
  "chd                                     ",
  "chd                                     ",
  "chd                                     ",
  "chd                                     " ;

 chd_0_iper = 1 ;
}
